`include "common.sv"
`include "asynch.v"
`include "wr_tx.sv"
`include "wr_gen.sv"
`include "fifo_intrf.sv"
`include "wr_bfm.sv"
`include "wr_mon.sv"
`include "wr_cov.sv"
`include "wr_agen.sv"
`include "rd_tx.sv"
`include "rd_gen.sv"
`include "rd_bfm.sv"
`include "rd_mon.sv"
`include "rd_cov.sv"
`include "rd_agent.sv"
`include "sbd.sv"
`include "env.sv"
`include "tb.sv"

